<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>5.0323,-7.75,102.993,-56.25</PageViewport>
<gate>
<ID>1</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>55,-52</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>4 </input>
<input>
<ID>IN_3</ID>5 </input>
<input>
<ID>IN_4</ID>6 </input>
<input>
<ID>IN_5</ID>7 </input>
<input>
<ID>IN_6</ID>7 </input>
<input>
<ID>IN_7</ID>7 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>2</ID>
<type>AE_FULLADDER_4BIT</type>
<position>40,-25</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>27 </input>
<input>
<ID>IN_2</ID>26 </input>
<input>
<ID>IN_3</ID>25 </input>
<input>
<ID>IN_B_0</ID>34 </input>
<input>
<ID>IN_B_1</ID>31 </input>
<input>
<ID>IN_B_2</ID>30 </input>
<input>
<ID>IN_B_3</ID>29 </input>
<output>
<ID>OUT_0</ID>1 </output>
<output>
<ID>OUT_1</ID>20 </output>
<output>
<ID>OUT_2</ID>21 </output>
<output>
<ID>OUT_3</ID>22 </output>
<input>
<ID>carry_in</ID>17 </input>
<output>
<ID>carry_out</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>3</ID>
<type>FF_GND</type>
<position>45,-50</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>23.5,-42.5</position>
<gparam>LABEL_TEXT Binary</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>77.5,-34</position>
<gparam>LABEL_TEXT Decimal</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>55,-44.5</position>
<gparam>LABEL_TEXT Hexadecimal</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>FF_GND</type>
<position>50,-27</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>29,-43</position>
<input>
<ID>N_in2</ID>6 </input>
<input>
<ID>N_in3</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>32,-43</position>
<input>
<ID>N_in2</ID>5 </input>
<input>
<ID>N_in3</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>35,-43</position>
<input>
<ID>N_in2</ID>4 </input>
<input>
<ID>N_in3</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>38,-43</position>
<input>
<ID>N_in2</ID>3 </input>
<input>
<ID>N_in3</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>41,-43</position>
<input>
<ID>N_in2</ID>2 </input>
<input>
<ID>N_in3</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>32,-12</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>32,-18</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>39,-15</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>32,-15</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>39,-12</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>39,-18</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>32,-9</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>39,-9</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>27,-8.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>27,-11.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>27,-14.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>27,-17.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>47,-8.5</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>47,-11.5</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>47,-14.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>47,-17.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>78,-42</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>136 </input>
<input>
<ID>IN_2</ID>137 </input>
<input>
<ID>IN_3</ID>138 </input>
<input>
<ID>IN_4</ID>139 </input>
<input>
<ID>IN_5</ID>140 </input>
<input>
<ID>IN_6</ID>141 </input>
<input>
<ID>IN_7</ID>142 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>137</ID>
<type>AA_LABEL</type>
<position>29,-45</position>
<gparam>LABEL_TEXT S4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>32,-45</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>35,-45</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AA_LABEL</type>
<position>38,-45</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>AA_LABEL</type>
<position>41,-45</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>AE_RAM_8x8</type>
<position>62,-30</position>
<input>
<ID>ADDRESS_0</ID>1 </input>
<input>
<ID>ADDRESS_1</ID>20 </input>
<input>
<ID>ADDRESS_2</ID>21 </input>
<input>
<ID>ADDRESS_3</ID>22 </input>
<input>
<ID>ADDRESS_4</ID>23 </input>
<input>
<ID>ADDRESS_5</ID>146 </input>
<input>
<ID>ADDRESS_6</ID>146 </input>
<input>
<ID>ADDRESS_7</ID>146 </input>
<input>
<ID>DATA_IN_0</ID>135 </input>
<input>
<ID>DATA_IN_1</ID>136 </input>
<input>
<ID>DATA_IN_2</ID>137 </input>
<input>
<ID>DATA_IN_3</ID>138 </input>
<input>
<ID>DATA_IN_4</ID>139 </input>
<input>
<ID>DATA_IN_5</ID>140 </input>
<input>
<ID>DATA_IN_6</ID>141 </input>
<input>
<ID>DATA_IN_7</ID>142 </input>
<output>
<ID>DATA_OUT_0</ID>135 </output>
<output>
<ID>DATA_OUT_1</ID>136 </output>
<output>
<ID>DATA_OUT_2</ID>137 </output>
<output>
<ID>DATA_OUT_3</ID>138 </output>
<output>
<ID>DATA_OUT_4</ID>139 </output>
<output>
<ID>DATA_OUT_5</ID>140 </output>
<output>
<ID>DATA_OUT_6</ID>141 </output>
<output>
<ID>DATA_OUT_7</ID>142 </output>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:1 1</lparam>
<lparam>Address:2 2</lparam>
<lparam>Address:3 3</lparam>
<lparam>Address:4 4</lparam>
<lparam>Address:5 5</lparam>
<lparam>Address:6 6</lparam>
<lparam>Address:7 7</lparam>
<lparam>Address:8 8</lparam>
<lparam>Address:9 9</lparam>
<lparam>Address:10 16</lparam>
<lparam>Address:11 17</lparam>
<lparam>Address:12 18</lparam>
<lparam>Address:13 19</lparam>
<lparam>Address:14 20</lparam>
<lparam>Address:15 21</lparam>
<lparam>Address:16 22</lparam>
<lparam>Address:17 23</lparam>
<lparam>Address:18 24</lparam>
<lparam>Address:19 25</lparam>
<lparam>Address:20 32</lparam>
<lparam>Address:21 33</lparam>
<lparam>Address:22 34</lparam>
<lparam>Address:23 35</lparam>
<lparam>Address:24 36</lparam>
<lparam>Address:25 37</lparam>
<lparam>Address:26 38</lparam>
<lparam>Address:27 39</lparam>
<lparam>Address:28 40</lparam>
<lparam>Address:29 41</lparam>
<lparam>Address:30 48</lparam>
<lparam>Address:31 49</lparam></gate>
<gate>
<ID>144</ID>
<type>FF_GND</type>
<position>53.5,-28.5</position>
<output>
<ID>OUT_0</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-36,41.5,-29</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-36 2</intersection>
<intersection>-33.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>41,-42,41,-36</points>
<connection>
<GID>22</GID>
<name>N_in3</name></connection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>41,-36,41.5,-36</points>
<intersection>41 1</intersection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>41.5,-33.5,57,-33.5</points>
<connection>
<GID>143</GID>
<name>ADDRESS_0</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-55,41,-44</points>
<connection>
<GID>22</GID>
<name>N_in2</name></connection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-55,50,-55</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-54,38,-44</points>
<connection>
<GID>20</GID>
<name>N_in2</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-54,50,-54</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-53,35,-44</points>
<connection>
<GID>18</GID>
<name>N_in2</name></connection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-53,50,-53</points>
<connection>
<GID>1</GID>
<name>IN_2</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-52,32,-44</points>
<connection>
<GID>16</GID>
<name>N_in2</name></connection>
<intersection>-52 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-52,50,-52</points>
<connection>
<GID>1</GID>
<name>IN_3</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-51,29,-44</points>
<connection>
<GID>14</GID>
<name>N_in2</name></connection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-51,50,-51</points>
<connection>
<GID>1</GID>
<name>IN_4</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-49,50,-49</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>50 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>50,-50,50,-48</points>
<connection>
<GID>1</GID>
<name>IN_5</name></connection>
<connection>
<GID>1</GID>
<name>IN_6</name></connection>
<connection>
<GID>1</GID>
<name>IN_7</name></connection>
<intersection>-49 1</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-26,50,-24</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-24,50,-24</points>
<connection>
<GID>2</GID>
<name>carry_in</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-42,38,-35</points>
<connection>
<GID>20</GID>
<name>N_in3</name></connection>
<intersection>-35 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>40.5,-35,40.5,-29</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>-35 2</intersection>
<intersection>-32.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>38,-35,40.5,-35</points>
<intersection>38 0</intersection>
<intersection>40.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>40.5,-32.5,57,-32.5</points>
<connection>
<GID>143</GID>
<name>ADDRESS_1</name></connection>
<intersection>40.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-34,39.5,-29</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>-34 2</intersection>
<intersection>-31.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>35,-42,35,-34</points>
<connection>
<GID>18</GID>
<name>N_in3</name></connection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35,-34,39.5,-34</points>
<intersection>35 1</intersection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>39.5,-31.5,57,-31.5</points>
<connection>
<GID>143</GID>
<name>ADDRESS_2</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-42,32,-33</points>
<connection>
<GID>16</GID>
<name>N_in3</name></connection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32,-33,38.5,-33</points>
<intersection>32 0</intersection>
<intersection>38.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>38.5,-33,38.5,-29</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>-33 2</intersection>
<intersection>-30.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>38.5,-30.5,57,-30.5</points>
<connection>
<GID>143</GID>
<name>ADDRESS_3</name></connection>
<intersection>38.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-42,29,-31.5</points>
<connection>
<GID>14</GID>
<name>N_in3</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-31.5,31.5,-31.5</points>
<intersection>29 0</intersection>
<intersection>31.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>31.5,-31.5,31.5,-24</points>
<intersection>-31.5 1</intersection>
<intersection>-29.5 4</intersection>
<intersection>-24 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-24,32,-24</points>
<connection>
<GID>2</GID>
<name>carry_out</name></connection>
<intersection>31.5 2</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>31.5,-29.5,57,-29.5</points>
<connection>
<GID>143</GID>
<name>ADDRESS_4</name></connection>
<intersection>31.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-21,35,-9</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>-9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>34,-9,35,-9</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-21,36,-12</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-12,36,-12</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-21,37,-15</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-15,37,-15</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-21,38,-18</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-18,38,-18</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-21,42,-9</points>
<connection>
<GID>2</GID>
<name>IN_B_3</name></connection>
<intersection>-9 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>41,-9,42,-9</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-21,43,-12</points>
<connection>
<GID>2</GID>
<name>IN_B_2</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-12,43,-12</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-21,44,-15</points>
<connection>
<GID>2</GID>
<name>IN_B_1</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-15,44,-15</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-21,45,-18</points>
<connection>
<GID>2</GID>
<name>IN_B_0</name></connection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-18,45,-18</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-45,65.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_IN_0</name></connection>
<intersection>-45 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-45,73,-45</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65.5,-37,65.5,-37</points>
<intersection>65.5 0</intersection>
<intersection>65.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>65.5,-37,65.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-37 2</intersection></vsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-44,64.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_IN_1</name></connection>
<intersection>-44 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64.5,-44,73,-44</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-37,64.5,-37</points>
<intersection>64.5 0</intersection>
<intersection>64.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>64.5,-37,64.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-37 2</intersection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-43,63.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_IN_2</name></connection>
<intersection>-43 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-43,73,-43</points>
<connection>
<GID>53</GID>
<name>IN_2</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-37,63.5,-37</points>
<intersection>63.5 0</intersection>
<intersection>63.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>63.5,-37,63.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-37 2</intersection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-42,62.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_IN_3</name></connection>
<intersection>-42 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-42,73,-42</points>
<connection>
<GID>53</GID>
<name>IN_3</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-37,62.5,-37</points>
<intersection>62.5 0</intersection>
<intersection>62.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>62.5,-37,62.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-37 2</intersection></vsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61.5,-41,73,-41</points>
<connection>
<GID>53</GID>
<name>IN_4</name></connection>
<intersection>61.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>61.5,-41,61.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_IN_4</name></connection>
<intersection>-41 1</intersection>
<intersection>-37 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>61.5,-37,61.5,-37</points>
<intersection>61.5 5</intersection>
<intersection>61.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>61.5,-37,61.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_OUT_4</name></connection>
<intersection>-37 6</intersection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-40,60.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_IN_5</name></connection>
<intersection>-40 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-40,73,-40</points>
<connection>
<GID>53</GID>
<name>IN_5</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60.5,-37,60.5,-37</points>
<intersection>60.5 0</intersection>
<intersection>60.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>60.5,-37,60.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_OUT_5</name></connection>
<intersection>-37 2</intersection></vsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-39,59.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_IN_6</name></connection>
<intersection>-39 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-39,73,-39</points>
<connection>
<GID>53</GID>
<name>IN_6</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59.5,-37,59.5,-37</points>
<intersection>59.5 0</intersection>
<intersection>59.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>59.5,-37,59.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_OUT_6</name></connection>
<intersection>-37 2</intersection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-38,58.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_IN_7</name></connection>
<intersection>-38 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-38,73,-38</points>
<connection>
<GID>53</GID>
<name>IN_7</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>58.5,-37,58.5,-37</points>
<intersection>58.5 0</intersection>
<intersection>58.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>58.5,-37,58.5,-37</points>
<connection>
<GID>143</GID>
<name>DATA_OUT_7</name></connection>
<intersection>-37 2</intersection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-27.5,57,-27.5</points>
<connection>
<GID>144</GID>
<name>OUT_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-28.5,57,-26.5</points>
<intersection>-28.5 3</intersection>
<intersection>-27.5 1</intersection>
<intersection>-27.5 4</intersection>
<intersection>-26.5 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>57,-28.5,57,-28.5</points>
<connection>
<GID>143</GID>
<name>ADDRESS_5</name></connection>
<intersection>57 2</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>57,-27.5,57,-27.5</points>
<connection>
<GID>143</GID>
<name>ADDRESS_6</name></connection>
<intersection>57 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>57,-26.5,57,-26.5</points>
<connection>
<GID>143</GID>
<name>ADDRESS_7</name></connection>
<intersection>57 2</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,33.6692,338.954,-134.146</PageViewport></page 1>
<page 2>
<PageViewport>0,33.6692,338.954,-134.146</PageViewport></page 2>
<page 3>
<PageViewport>0,33.6692,338.954,-134.146</PageViewport></page 3>
<page 4>
<PageViewport>0,33.6692,338.954,-134.146</PageViewport></page 4>
<page 5>
<PageViewport>0,33.6692,338.954,-134.146</PageViewport></page 5>
<page 6>
<PageViewport>0,33.6692,338.954,-134.146</PageViewport></page 6>
<page 7>
<PageViewport>0,33.6692,338.954,-134.146</PageViewport></page 7>
<page 8>
<PageViewport>0,33.6692,338.954,-134.146</PageViewport></page 8>
<page 9>
<PageViewport>0,33.6692,338.954,-134.146</PageViewport></page 9></circuit>